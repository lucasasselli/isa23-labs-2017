package tta0_imem_mau is
   -- created by generatebits
   constant IMEMMAUWIDTH : positive := 84;
end tta0_imem_mau;
