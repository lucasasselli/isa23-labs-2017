package tta0_imem_mau is
   -- created by generatebits
   constant IMEMMAUWIDTH : positive := 42;
end tta0_imem_mau;
