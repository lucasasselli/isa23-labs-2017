package tta0_imem_mau is
   -- created by generatebits
   constant IMEMMAUWIDTH : positive := 126;
end tta0_imem_mau;
