package tta0_params is
  constant fu_LSU_dataw : integer := 32;
  constant fu_LSU_addrw : integer := 16;
end tta0_params;
